module Control (
    
);

endmodule
