module Processor(
    input clk  
);


endmodule
